-- hier steht unser System, an welches noch IO, Mem und clk, rst hinkommen (auch die TB)

ENtity System IS

END Entity;

Architecture behav of System IS

END Architecture;

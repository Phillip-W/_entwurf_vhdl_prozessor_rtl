-- Hier wird die Verkabelung der einzlnen Komponenten statt finden, aber keine eigene Logik!
